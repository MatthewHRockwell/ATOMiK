// =============================================================================
// ATOMiK Delta Accumulator Module
// 
// Module:      atomik_delta_acc
// Description: Maintains initial state and accumulates deltas via XOR composition
// 
// Key Features:
//   - Dual-register architecture (initial_state, delta_accumulator)
//   - Single-cycle XOR accumulation (no carry propagation)
//   - Configurable delta width (64-bit default)
//   - Synchronous reset to known state
//   - Zero detection for delta algebra verification
//
// Mathematical Foundation (from Phase 1 Lean4 proofs):
//   - delta_comm:        δ₁ ⊕ δ₂ = δ₂ ⊕ δ₁ (order irrelevant)
//   - delta_assoc:       (δ₁ ⊕ δ₂) ⊕ δ₃ = δ₁ ⊕ (δ₂ ⊕ δ₃) (grouping irrelevant)
//   - delta_self_inverse: δ ⊕ δ = 0 (enables undo/verification)
//
// Performance:
//   - Accumulate latency: 1 clock cycle
//   - Load latency: 1 clock cycle
//   - Throughput: 1 delta per cycle (back-to-back supported)
//
// Target: Gowin GW1NR-9 (Tang Nano 9K)
// Author: ATOMiK Project
// Date:   January 25, 2026
// =============================================================================

`timescale 1ns / 1ps

module atomik_delta_acc #(
    parameter DELTA_WIDTH = 64      // Width of delta and state (matches Phase 1 proofs)
)(
    // Clock and Reset
    input  wire                     clk,            // System clock
    input  wire                     rst_n,          // Active-low synchronous reset
    
    // Delta Input Interface
    input  wire [DELTA_WIDTH-1:0]   delta_in,       // Delta value to accumulate
    input  wire                     delta_valid,    // Delta input valid strobe
    
    // Initial State Interface
    input  wire [DELTA_WIDTH-1:0]   initial_state_in,   // New initial state value
    input  wire                     load_initial,       // Load initial state strobe
    
    // Output Interface
    output wire [DELTA_WIDTH-1:0]   initial_state_out,      // Current initial state
    output wire [DELTA_WIDTH-1:0]   delta_accumulator_out,  // Current accumulated delta
    
    // Status Interface
    output wire                     accumulator_zero    // High when accumulator = 0
);

    // =========================================================================
    // Internal Registers
    // =========================================================================
    
    // Initial state register: S₀ from which all deltas are applied
    // Updated only on LOAD operation
    reg [DELTA_WIDTH-1:0] initial_state;
    
    // Delta accumulator: Running XOR composition of all deltas
    // δ_acc = δ₁ ⊕ δ₂ ⊕ ... ⊕ δₙ
    // Updated on each ACCUMULATE operation
    reg [DELTA_WIDTH-1:0] delta_accumulator;

    // =========================================================================
    // Main Sequential Logic
    // =========================================================================
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            // Synchronous reset: Clear both registers
            // This establishes a known starting state
            initial_state     <= {DELTA_WIDTH{1'b0}};
            delta_accumulator <= {DELTA_WIDTH{1'b0}};
        end
        else begin
            // Load initial state - also clears delta accumulator
            // This establishes a fresh starting point
            if (load_initial) begin
                initial_state     <= initial_state_in;
                delta_accumulator <= {DELTA_WIDTH{1'b0}};  // Clear accumulator on LOAD
            end
            
            // Accumulate delta via XOR
            // Key insight: XOR has no carry propagation, so this is
            // a single-cycle operation even for 64-bit width
            if (delta_valid) begin
                delta_accumulator <= delta_accumulator ^ delta_in;
            end
        end
    end

    // =========================================================================
    // Output Assignments
    // =========================================================================
    
    // Direct register outputs
    assign initial_state_out     = initial_state;
    assign delta_accumulator_out = delta_accumulator;
    
    // Zero detection: OR-reduction followed by inversion
    // This implements the check for δ_acc = 0, which is useful for:
    //   1. Verifying δ ⊕ δ = 0 (self-inverse property)
    //   2. Detecting when state equals initial_state
    //   3. Debugging and verification
    //
    // Implementation: ~(|delta_accumulator) is a tree of OR gates
    // followed by an inverter, typically ~8 LUTs for 64-bit input
    assign accumulator_zero = ~(|delta_accumulator);

    // =========================================================================
    // Assertions (for simulation only)
    // =========================================================================
    
    `ifdef SIMULATION
    // Verify self-inverse property: accumulating same delta twice should
    // return accumulator to previous state
    reg [DELTA_WIDTH-1:0] prev_accumulator;
    reg [DELTA_WIDTH-1:0] prev_delta;
    reg                   check_self_inverse;
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            prev_accumulator   <= {DELTA_WIDTH{1'b0}};
            prev_delta         <= {DELTA_WIDTH{1'b0}};
            check_self_inverse <= 1'b0;
        end
        else if (delta_valid) begin
            prev_accumulator <= delta_accumulator;
            prev_delta       <= delta_in;
            
            // Check if this delta equals the previous one
            if (delta_in == prev_delta && check_self_inverse) begin
                // After δ ⊕ δ, accumulator should equal prev_accumulator
                // (two applications of same delta cancel out)
                // Note: This check happens one cycle late, which is correct
            end
            check_self_inverse <= 1'b1;
        end
    end
    `endif

endmodule

// =============================================================================
// Module Documentation
// =============================================================================
//
// USAGE EXAMPLE:
// --------------
// atomik_delta_acc #(
//     .DELTA_WIDTH(64)
// ) u_delta_acc (
//     .clk                 (clk),
//     .rst_n               (rst_n),
//     .delta_in            (delta_value),
//     .delta_valid         (delta_strobe),
//     .initial_state_in    (new_initial_state),
//     .load_initial        (load_strobe),
//     .initial_state_out   (current_initial),
//     .delta_accumulator_out(current_accumulator),
//     .accumulator_zero    (acc_is_zero)
// );
//
// TIMING DIAGRAMS:
// ----------------
// Load Operation:
//   clk:          __|‾‾|__|‾‾|__|‾‾|__
//   load_initial: __|‾‾‾‾‾|________
//   initial_in:   XX|INIT |XXXXXXXX
//   initial_out:  00|0000 |INIT----
//
// Accumulate Operation:
//   clk:          __|‾‾|__|‾‾|__|‾‾|__
//   delta_valid:  __|‾‾‾‾‾|‾‾‾‾‾|____
//   delta_in:     XX| δ1  | δ2  |XXXX
//   accum_out:    00| δ1  |δ1⊕δ2|----
//
// RESOURCE ESTIMATES (GW1NR-9):
// -----------------------------
//   Flip-Flops: 128 (64 + 64)
//   LUTs:       ~82 (64 XOR + 10 control + 8 zero detect)
//   Fmax:       >300 MHz (XOR has no carry chain)
//
// =============================================================================
